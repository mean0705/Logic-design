library verilog;
use verilog.vl_types.all;
entity Total is
end Total;
